write back a file or signal
